module abs

pub fn add_m(x int, y int) int {
	return x + y
}
