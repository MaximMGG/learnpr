module main

import abs

fn main() {
	println('Main module')
	println(abs.add_m(1, 2))
}
